`timescale 1ns / 1 ps
module (   // translated from Lola
endmodule
